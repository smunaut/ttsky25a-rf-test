MACRO tt_um_tnt_rf_test
  CLASS BLOCK ;
  FOREIGN tt_um_tnt_rf_test ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.000 10.000 23.000 217.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.000 10.000 43.000 217.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.000 10.000 63.000 217.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.000 10.000 127.000 217.500 ;
    END
  END VGND
  PIN VDPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 25.000 10.000 27.000 217.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.000 10.000 47.000 217.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 65.000 10.000 67.000 217.500 ;
    END
  END VDPWR
  PIN VDPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 129.000 10.000 131.000 217.500 ;
    END
  END VDPWR
  OBS
      LAYER nwell ;
        RECT 6.165 35.000 154.835 223.305 ;
      LAYER li1 ;
        RECT 6.165 35.190 154.835 223.115 ;
      LAYER met1 ;
        RECT 6.010 35.190 154.990 223.115 ;
      LAYER met2 ;
        RECT 6.010 37.130 154.990 224.735 ;
      LAYER met3 ;
        RECT 6.010 56.440 154.990 224.800 ;
      LAYER met4 ;
        RECT 18.440 224.360 30.270 224.775 ;
        RECT 31.370 224.360 33.030 224.775 ;
        RECT 34.130 224.360 35.790 224.775 ;
        RECT 36.890 224.360 38.550 224.775 ;
        RECT 39.650 224.360 41.310 224.775 ;
        RECT 42.410 224.360 44.070 224.775 ;
        RECT 45.170 224.360 46.830 224.775 ;
        RECT 47.930 224.360 49.590 224.775 ;
        RECT 50.690 224.360 52.350 224.775 ;
        RECT 53.450 224.360 55.110 224.775 ;
        RECT 56.210 224.360 57.870 224.775 ;
        RECT 58.970 224.360 60.630 224.775 ;
        RECT 61.730 224.360 63.390 224.775 ;
        RECT 64.490 224.360 66.150 224.775 ;
        RECT 67.250 224.360 68.910 224.775 ;
        RECT 70.010 224.360 71.670 224.775 ;
        RECT 72.770 224.360 74.430 224.775 ;
        RECT 75.530 224.360 77.190 224.775 ;
        RECT 78.290 224.360 79.950 224.775 ;
        RECT 81.050 224.360 82.710 224.775 ;
        RECT 83.810 224.360 85.470 224.775 ;
        RECT 86.570 224.360 88.230 224.775 ;
        RECT 89.330 224.360 90.990 224.775 ;
        RECT 92.090 224.360 93.750 224.775 ;
        RECT 94.850 224.360 96.510 224.775 ;
        RECT 97.610 224.360 99.270 224.775 ;
        RECT 100.370 224.360 102.030 224.775 ;
        RECT 103.130 224.360 104.790 224.775 ;
        RECT 105.890 224.360 107.550 224.775 ;
        RECT 108.650 224.360 110.310 224.775 ;
        RECT 111.410 224.360 113.070 224.775 ;
        RECT 114.170 224.360 115.830 224.775 ;
        RECT 116.930 224.360 118.590 224.775 ;
        RECT 119.690 224.360 121.350 224.775 ;
        RECT 122.450 224.360 124.110 224.775 ;
        RECT 125.210 224.360 126.870 224.775 ;
        RECT 127.970 224.360 129.630 224.775 ;
        RECT 130.730 224.360 132.390 224.775 ;
        RECT 133.490 224.360 135.150 224.775 ;
        RECT 136.250 224.360 137.910 224.775 ;
        RECT 139.010 224.360 140.670 224.775 ;
        RECT 141.770 224.360 143.430 224.775 ;
        RECT 144.530 224.360 146.190 224.775 ;
        RECT 147.290 224.360 150.865 224.775 ;
        RECT 18.440 217.900 150.865 224.360 ;
        RECT 18.440 77.335 20.600 217.900 ;
        RECT 23.400 77.335 24.600 217.900 ;
        RECT 27.400 77.335 40.600 217.900 ;
        RECT 43.400 77.335 44.600 217.900 ;
        RECT 47.400 77.335 60.600 217.900 ;
        RECT 63.400 77.335 64.600 217.900 ;
        RECT 67.400 77.335 124.600 217.900 ;
        RECT 127.400 77.335 128.600 217.900 ;
        RECT 131.400 77.335 150.865 217.900 ;
  END
END tt_um_tnt_rf_test
END LIBRARY

